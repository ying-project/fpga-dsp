// Original VHDL source code Copyright 1995-2021 DOULOS
// Modified by: Zhiying Meng